`ifndef MOBILENET_DEFINES_VH
`define MOBILENET_DEFINES_VH

// ============================================================
// MobileNetV1 ȫ�ֲ������� (32��32 PE����)
// ============================================================

// -------------------- ����λ�� --------------------
`define DATA_W      8      // INT8
`define ACC_W       32     // �ۼ���λ��
`define WEIGHT_W    8      // Ȩ��λ��
`define PSUM_W      18     // ���ֺ�λ��
`define PROD_W      16     // �˻�λ��

// -------------------- PE�������� (32��32) --------------------
`define PE_ROWS     32
`define PE_COLS     32
`define UNIT_NUM    32
`define LANES       32

// -------------------- MobileNetV1 ������ --------------------
`define TOTAL_LAYERS              29     // Layer 0-28 (��29��)
`define MAX_LAYER_ID              28
`define TOTAL_CONV_DW_PW_LAYERS   27

// -------------------- ͼ��ߴ����� --------------------
`define MAX_IMG_W     224
`define MAX_IMG_H     224
`define MAX_CHANNELS  1024
`define MAX_OUT_W     112
`define MAX_OUT_H     112

// -------------------- ����ͼ��������� --------------------
// (112*112*64 / 16 = 50176 words)
`define FEATURE_BUF_DEPTH  50176

// -------------------- Ȩ�ش洢����ַ --------------------
`define L0_WEIGHT_BASE   9'd0     // Layer0 �� 0 ��ʼ
`define L2_WEIGHT_BASE   9'd64    // Layer2 �� 64 ��ʼ

// -------------------- ����·�� --------------------
`define DATA_PATH  "D:/NoC/mycode/mobilenet_acc2/data/"

// ============================================================
// Layer Type Definitions (3-bit)
// ============================================================
`define LAYER_TYPE_CONV   3'd0    // ��һ����׼3x3���
`define LAYER_TYPE_DW     3'd1    // Depthwise Convolution
`define LAYER_TYPE_PW     3'd2    // Pointwise Convolution
`define LAYER_TYPE_AP     3'd3    // Global Average Pooling
`define LAYER_TYPE_FC     3'd4    // Fully Connected

// ============================================================
// Memory Parameters
// ============================================================
`define WEIGHT_ADDR_W   16
`define BIAS_ADDR_W     12
`define FEAT_ADDR_W     17

// ============================================================
// Fast Simulation Parameters
// ============================================================
`define FAST_SIM_ENABLE  0    // Ĭ�Ϲر�
`define FAST_SIM_NO_MAC  0    // Ĭ�Ϲر�

`endif  // MOBILENET_DEFINES_VH
