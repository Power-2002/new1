`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/12/15 16:37:49
// Design Name: 
// Module Name: simple_column_scanner_pipeline
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module simple_column_scanner_pipeline #(
  parameter integer OUT_W   = 112,
  parameter integer OUT_H   = 112,
  parameter integer TILE_H  = 6,
  parameter integer K       = 3,
  parameter integer PADDING = 1  // ? �Ļ� 1����˫����һ�£�
)(
  input  wire clk,
  input  wire rst_n,
  input  wire start,

  // Runtime configuration
  input  wire [7:0] cfg_w,
  input  wire [7:0] cfg_h,
  input  wire       stride2_en,

  // ? �ָ���Щ�˿ڣ�������ı䣩
  output reg  [$clog2(OUT_H)-1:0] current_tile_row,  // ��ǰ tile ��
  output reg  tile_start,  // �� tile ��ʼ����
  input  wire buffer_ready,

  // Read interface
  output wire read_enable,
  output wire [$clog2(OUT_W)-1:0] read_addr,

  // Status
  output reg  busy,
  output reg  done,
  output reg  [$clog2(OUT_W)-1:0] current_col
);

  // ============================================================
  // ��������
  // ============================================================
  localparam integer STEP_ROW_S1_INT = (TILE_H - K + 1);      // 4
  localparam integer STEP_ROW_S2_INT = (TILE_H - K + 1) * 2;  // 8
  
  wire [$clog2(OUT_H)-1:0] step_row_s1 = STEP_ROW_S1_INT[$clog2(OUT_H)-1:0];
  wire [$clog2(OUT_H)-1:0] step_row_s2 = STEP_ROW_S2_INT[$clog2(OUT_H)-1:0];

  // ============================================================
  // ״̬�������� 2 ��״̬��
  // ============================================================
  localparam S_IDLE = 1'b0;
  localparam S_SCAN = 1'b1;

  reg state;
  reg [$clog2(OUT_W)-1:0] col_counter;

  // ============================================================
  // Runtime configuration
  // ============================================================
  wire [7:0] cfg_w_clamped = (cfg_w > OUT_W[7:0]) ? OUT_W[7:0] : cfg_w;
  wire [7:0] cfg_h_clamped = (cfg_h > OUT_H[7:0]) ? OUT_H[7:0] : cfg_h;

  // Padded width
  wire [$clog2(OUT_W)-1:0] padded_w = cfg_w_clamped[$clog2(OUT_W)-1:0] + (PADDING * 2);
  wire [$clog2(OUT_W)-1:0] w_minus1 = padded_w - 1'b1;
  wire [$clog2(OUT_W)-1:0] w_minus2 = (padded_w >= 2) ? (padded_w - 2'd2) : {($clog2(OUT_W)){1'b0}};
  
  wire [$clog2(OUT_H)-1:0] h_limit = cfg_h_clamped[$clog2(OUT_H)-1:0];

// ? ��ǰԤȡ�����㣨80% λ�ã�Ԥ�� 20% �ص�ʱ�䣩
wire [$clog2(OUT_W)-1:0] prefetch_trigger_col;
assign prefetch_trigger_col = (padded_w * 4) / 5;  // 80% λ��

// ? ����Ƿ�Ӧ����ǰԤȡ��һ�� tile
wire should_trigger_prefetch_s1 = (col_counter == prefetch_trigger_col) && 
                                   ((current_tile_row + step_row_s1) < h_limit) && 
                                   (! stride2_en);

wire should_trigger_prefetch_s2 = (col_counter == prefetch_trigger_col) && 
                                   ((current_tile_row + step_row_s2) < h_limit) && 
                                   (stride2_en);

  // ============================================================
  // Output assignments
  // ============================================================
  assign read_enable = (state == S_SCAN) && buffer_ready;
  assign read_addr   = col_counter;

  // ============================================================
  // ? �ؼ�������FSM ���� tile ����
  // ============================================================
  always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      state            <= S_IDLE;
      busy             <= 1'b0;
      done             <= 1'b0;
      col_counter      <= {($clog2(OUT_W)){1'b0}};
      current_col      <= {($clog2(OUT_W)){1'b0}};
      current_tile_row <= {($clog2(OUT_H)){1'b0}};
      tile_start       <= 1'b0;
    end else begin
      done       <= 1'b0;  // Pulse
      tile_start <= 1'b0;  // Pulse

      case (state)
        
        // ========================================
        // IDLE: Wait for start
        // ========================================
        S_IDLE: begin
          busy             <= 1'b0;
          col_counter      <= 0;
          current_col      <= 0;
          current_tile_row <= 0;

          if (start) begin
            busy       <= 1'b1;
            tile_start <= 1'b1;  // ? ������һ�� tile Ԥȡ
            state      <= S_SCAN;
          end
        end

        // ========================================
        // SCAN: Scan columns with tile iteration
        // ========================================
// ========== �滻�� 106-156 �е� S_SCAN ״̬�� ==========

S_SCAN: begin
  if (buffer_ready) begin
    current_col <= col_counter;

    // ? ��ǰԤȡ�߼�����ɨ�赽 80% ʱ�ʹ�����һ�� tile ��Ԥȡ
    if (should_trigger_prefetch_s1 || should_trigger_prefetch_s2) begin
      tile_start <= 1'b1;  // ? ��ǰ 20% �Ϳ�ʼԤȡ
    end

    // Stride = 1
    if (! stride2_en) begin
      if (col_counter < w_minus1) begin
        col_counter <= col_counter + 1'b1;
      end else begin
        // һ��ɨ����ɣ����� tile_row
        col_counter <= 0;
        
        if ((current_tile_row + step_row_s1) < h_limit) begin
          current_tile_row <= current_tile_row + step_row_s1;
          // ? ע�⣺���������ﴥ�� tile_start������ 80% ʱ��ǰ������
        end else begin
          // ���� tile ���
          busy  <= 1'b0;
          done  <= 1'b1;
          state <= S_IDLE;
        end
      end
    end
    
    // Stride = 2
    else begin
      if (col_counter < w_minus2) begin
        col_counter <= col_counter + 2'd2;
      end else begin
        col_counter <= 0;
        
        if ((current_tile_row + step_row_s2) < h_limit) begin
          current_tile_row <= current_tile_row + step_row_s2;
          // ? ���������ﴥ�� tile_start
        end else begin
          busy  <= 1'b0;
          done  <= 1'b1;
          state <= S_IDLE;
        end
      end
    end
  end
end

        default: state <= S_IDLE;
      endcase
    end
  end

endmodule